module plru;

endmodule