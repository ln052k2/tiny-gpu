// Logger class to help with testing

// Generates a log file with date/time stamp
// Appends to log file and displays messages to console