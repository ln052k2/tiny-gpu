// Uses helper module Memory -- similar to top module of a testbench

// Generate clock with a period of 25 us
// Reset DUT - wait one posedge of clock

// Load program and data memory

// Write number of threads to register device_control_data

// Start DUT and wait for it to finish