module plru;
endmodule