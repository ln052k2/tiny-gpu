  module memif_connector (
    mem_if.consumer consumer_if,
    mem_if.mem memory_if 
);