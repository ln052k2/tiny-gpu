package alu_state_pkg;
    typedef enum logic [1:0] {IDLE, WAIT_DIV, DONE} alu_state_t;
endpackage