// Program memory: 8 address bits, 16 data bits, 1 channel
// TODO: Move program instruction sequence to separate file (?)

// Data memory: 8 address bits, 8 data bits, 4 channels
// Matrix A and B are both [0, 1, 2, 3, 4, 5, 6, 7]

// 8 threads